library verilog;
use verilog.vl_types.all;
entity Controlsalida_tiempos_tb is
end Controlsalida_tiempos_tb;
