library verilog;
use verilog.vl_types.all;
entity empaquetado is
end empaquetado;
